library verilog;
use verilog.vl_types.all;
entity Absl_vlg_vec_tst is
end Absl_vlg_vec_tst;
