library verilog;
use verilog.vl_types.all;
entity IndexRegister_vlg_vec_tst is
end IndexRegister_vlg_vec_tst;
