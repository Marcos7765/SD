library verilog;
use verilog.vl_types.all;
entity SAD_vlg_vec_tst is
end SAD_vlg_vec_tst;
