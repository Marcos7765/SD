library verilog;
use verilog.vl_types.all;
entity CustomAdder_vlg_vec_tst is
end CustomAdder_vlg_vec_tst;
