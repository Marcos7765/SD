library verilog;
use verilog.vl_types.all;
entity DataRegister_vlg_vec_tst is
end DataRegister_vlg_vec_tst;
