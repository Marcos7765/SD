library verilog;
use verilog.vl_types.all;
entity CustomAdder_vlg_check_tst is
    port(
        Result          : in     vl_logic_vector(31 downto 0);
        sampler_rx      : in     vl_logic
    );
end CustomAdder_vlg_check_tst;
