library verilog;
use verilog.vl_types.all;
entity Comparator_vlg_check_tst is
    port(
        Output          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Comparator_vlg_check_tst;
