LIBRARY ieee;
USE ieee.std_logic_1164.all;
--diretamente do velho lab de cd
ENTITY decod7seg IS
PORT(
	A: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	S : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END;
ARCHITECTURE main OF decod7seg IS
BEGIN
	WITH A SELECT
		S <= "1000000" WHEN "0000",
			"1111001" WHEN "0001",
			"0100100" WHEN "0010",
			"0110000" WHEN "0011",
			"0011001" WHEN "0100",
			"0010010" WHEN "0101",
			"0000010" WHEN "0110",
			"1111000" WHEN "0111",
			"0000000" WHEN "1000",
			"0010000" WHEN "1001",
			"1111111" WHEN OTHERS;
END;